module uart_macro_wrapper (
`ifdef USE_POWER_PINS
    inout vccd1,    // User area 1 1.8V supply
    inout vssd1,    // User area 1 digital ground
`endif

    // Wishbone Slave ports
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // UART pins
    input uart_rx,
    output uart_tx,
    output [1:0] io_oeb,
    
    // IRQ
    output uart_irq
);

    // Instantiate CF_UART with Wishbone interface
    CF_UART_WB uart (
        .clk_i(wb_clk_i),
        .rst_i(wb_rst_i),
        .adr_i(wbs_adr_i),
        .dat_i(wbs_dat_i),
        .dat_o(wbs_dat_o),
        .sel_i(wbs_sel_i),
        .cyc_i(wbs_cyc_i),
        .stb_i(wbs_stb_i),
        .ack_o(wbs_ack_o),
        .we_i(wbs_we_i),
        .IRQ(uart_irq),
        .rx(uart_rx),
        .tx(uart_tx)
    );

    assign io_oeb[0] = 1'b1;
    assign io_oeb[1] = 1'b0;

endmodule